-------------------------------------------------------------------------------
-- system_my_peripheral_lab4_0_wrapper.vhd
-------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

library my_peripheral_lab4_v1_00_a;
use my_peripheral_lab4_v1_00_a.all;

entity system_my_peripheral_lab4_0_wrapper is
  port (
    S_AXI_ACLK : in std_logic;
    S_AXI_ARESETN : in std_logic;
    S_AXI_AWADDR : in std_logic_vector(31 downto 0);
    S_AXI_AWVALID : in std_logic;
    S_AXI_WDATA : in std_logic_vector(31 downto 0);
    S_AXI_WSTRB : in std_logic_vector(3 downto 0);
    S_AXI_WVALID : in std_logic;
    S_AXI_BREADY : in std_logic;
    S_AXI_ARADDR : in std_logic_vector(31 downto 0);
    S_AXI_ARVALID : in std_logic;
    S_AXI_RREADY : in std_logic;
    S_AXI_ARREADY : out std_logic;
    S_AXI_RDATA : out std_logic_vector(31 downto 0);
    S_AXI_RRESP : out std_logic_vector(1 downto 0);
    S_AXI_RVALID : out std_logic;
    S_AXI_WREADY : out std_logic;
    S_AXI_BRESP : out std_logic_vector(1 downto 0);
    S_AXI_BVALID : out std_logic;
    S_AXI_AWREADY : out std_logic;
    CLK_I : in std_logic;
    RESET_N_I : in std_logic;
    DIRECT_MODE_I : in std_logic;
    DISPLAY_MODE_I : in std_logic_vector(1 downto 0);
    VGA_HSYNC_O : out std_logic;
    VGA_VSYNC_O : out std_logic;
    BLANK_O : out std_logic;
    PIX_CLOCK_O : out std_logic;
    PSAVE_O : out std_logic;
    SYNC_O : out std_logic;
    RED_O : out std_logic_vector(7 downto 0);
    GREEN_O : out std_logic_vector(7 downto 0);
    BLUE_O : out std_logic_vector(7 downto 0)
  );
end system_my_peripheral_lab4_0_wrapper;

architecture STRUCTURE of system_my_peripheral_lab4_0_wrapper is

  component my_peripheral_lab4 is
    generic (
      C_S_AXI_DATA_WIDTH : INTEGER;
      C_S_AXI_ADDR_WIDTH : INTEGER;
      C_S_AXI_MIN_SIZE : std_logic_vector;
      C_USE_WSTRB : INTEGER;
      C_DPHASE_TIMEOUT : INTEGER;
      C_BASEADDR : std_logic_vector;
      C_HIGHADDR : std_logic_vector;
      C_FAMILY : STRING;
      C_NUM_REG : INTEGER;
      C_NUM_MEM : INTEGER;
      C_SLV_AWIDTH : INTEGER;
      C_SLV_DWIDTH : INTEGER
    );
    port (
      S_AXI_ACLK : in std_logic;
      S_AXI_ARESETN : in std_logic;
      S_AXI_AWADDR : in std_logic_vector((C_S_AXI_ADDR_WIDTH-1) downto 0);
      S_AXI_AWVALID : in std_logic;
      S_AXI_WDATA : in std_logic_vector((C_S_AXI_DATA_WIDTH-1) downto 0);
      S_AXI_WSTRB : in std_logic_vector(((C_S_AXI_DATA_WIDTH/8)-1) downto 0);
      S_AXI_WVALID : in std_logic;
      S_AXI_BREADY : in std_logic;
      S_AXI_ARADDR : in std_logic_vector((C_S_AXI_ADDR_WIDTH-1) downto 0);
      S_AXI_ARVALID : in std_logic;
      S_AXI_RREADY : in std_logic;
      S_AXI_ARREADY : out std_logic;
      S_AXI_RDATA : out std_logic_vector((C_S_AXI_DATA_WIDTH-1) downto 0);
      S_AXI_RRESP : out std_logic_vector(1 downto 0);
      S_AXI_RVALID : out std_logic;
      S_AXI_WREADY : out std_logic;
      S_AXI_BRESP : out std_logic_vector(1 downto 0);
      S_AXI_BVALID : out std_logic;
      S_AXI_AWREADY : out std_logic;
      CLK_I : in std_logic;
      RESET_N_I : in std_logic;
      DIRECT_MODE_I : in std_logic;
      DISPLAY_MODE_I : in std_logic_vector(1  downto  0);
      VGA_HSYNC_O : out std_logic;
      VGA_VSYNC_O : out std_logic;
      BLANK_O : out std_logic;
      PIX_CLOCK_O : out std_logic;
      PSAVE_O : out std_logic;
      SYNC_O : out std_logic;
      RED_O : out std_logic_vector(7  downto  0);
      GREEN_O : out std_logic_vector(7  downto  0);
      BLUE_O : out std_logic_vector(7  downto  0)
    );
  end component;

begin

  my_peripheral_lab4_0 : my_peripheral_lab4
    generic map (
      C_S_AXI_DATA_WIDTH => 32,
      C_S_AXI_ADDR_WIDTH => 32,
      C_S_AXI_MIN_SIZE => X"000001ff",
      C_USE_WSTRB => 0,
      C_DPHASE_TIMEOUT => 8,
      C_BASEADDR => X"7b200000",
      C_HIGHADDR => X"7b20ffff",
      C_FAMILY => "spartan6",
      C_NUM_REG => 1,
      C_NUM_MEM => 1,
      C_SLV_AWIDTH => 32,
      C_SLV_DWIDTH => 32
    )
    port map (
      S_AXI_ACLK => S_AXI_ACLK,
      S_AXI_ARESETN => S_AXI_ARESETN,
      S_AXI_AWADDR => S_AXI_AWADDR,
      S_AXI_AWVALID => S_AXI_AWVALID,
      S_AXI_WDATA => S_AXI_WDATA,
      S_AXI_WSTRB => S_AXI_WSTRB,
      S_AXI_WVALID => S_AXI_WVALID,
      S_AXI_BREADY => S_AXI_BREADY,
      S_AXI_ARADDR => S_AXI_ARADDR,
      S_AXI_ARVALID => S_AXI_ARVALID,
      S_AXI_RREADY => S_AXI_RREADY,
      S_AXI_ARREADY => S_AXI_ARREADY,
      S_AXI_RDATA => S_AXI_RDATA,
      S_AXI_RRESP => S_AXI_RRESP,
      S_AXI_RVALID => S_AXI_RVALID,
      S_AXI_WREADY => S_AXI_WREADY,
      S_AXI_BRESP => S_AXI_BRESP,
      S_AXI_BVALID => S_AXI_BVALID,
      S_AXI_AWREADY => S_AXI_AWREADY,
      CLK_I => CLK_I,
      RESET_N_I => RESET_N_I,
      DIRECT_MODE_I => DIRECT_MODE_I,
      DISPLAY_MODE_I => DISPLAY_MODE_I,
      VGA_HSYNC_O => VGA_HSYNC_O,
      VGA_VSYNC_O => VGA_VSYNC_O,
      BLANK_O => BLANK_O,
      PIX_CLOCK_O => PIX_CLOCK_O,
      PSAVE_O => PSAVE_O,
      SYNC_O => SYNC_O,
      RED_O => RED_O,
      GREEN_O => GREEN_O,
      BLUE_O => BLUE_O
    );

end architecture STRUCTURE;

